LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY CPU_tb IS
END CPU_tb;

ARCHITECTURE test OF CPU_tb IS
  COMPONENT CPU
    PORT (
      CLOCK_50 : IN STD_LOGIC := '0';
      PONTO_OPERACAO : IN STD_LOGIC := '0';
      PONTO_ESCREVE_C : IN STD_LOGIC := '0';
      PONTO_HAB_WRITE : IN STD_LOGIC := '0';
      PONTO_HAB_READ : IN STD_LOGIC := '0';
      PONTO_HAB_RAM : IN STD_LOGIC := '0';
      PONTO_MUX_RT_IMEDIATO : IN STD_LOGIC := '0';
      PONTO_BEQ : IN STD_LOGIC := '0';
      PONTO_MUX_RT_RD : IN STD_LOGIC := '0';
      PONTO_MUX_ALU_RAM : IN STD_LOGIC := '0';
      PONTO_MUX_JMP : IN STD_LOGIC := '0'
    );
  END COMPONENT;

  SIGNAL W_CLK : STD_LOGIC := '0';
  SIGNAL W_PONTO_OPERACAO : STD_LOGIC := '0';
  SIGNAL W_PONTO_ESCREVE_C : STD_LOGIC := '0';
  SIGNAL W_PONTO_HAB_WRITE : STD_LOGIC := '0';
  SIGNAL W_PONTO_HAB_READ : STD_LOGIC := '0';
  SIGNAL W_PONTO_HAB_RAM : STD_LOGIC := '0';
  SIGNAL W_PONTO_MUX_RT_IMEDIATO : STD_LOGIC := '0';
  SIGNAL W_PONTO_BEQ : STD_LOGIC := '0';
  SIGNAL W_PONTO_MUX_RT_RD : STD_LOGIC := '0';
  SIGNAL W_PONTO_MUX_ALU_RAM : STD_LOGIC := '0';
  SIGNAL W_PONTO_MUX_JMP : STD_LOGIC := '0';

  CONSTANT PERIODO : TIME := 10 ps;

BEGIN

  TL : CPU
  PORT MAP(
    CLOCK_50 => W_CLK,
    PONTO_OPERACAO => W_PONTO_OPERACAO,
    PONTO_ESCREVE_C => W_PONTO_ESCREVE_C,
    PONTO_HAB_WRITE => W_PONTO_HAB_WRITE,
    PONTO_HAB_READ => W_PONTO_HAB_READ,
    PONTO_HAB_RAM => W_PONTO_HAB_RAM,
    PONTO_MUX_RT_IMEDIATO => W_PONTO_MUX_RT_IMEDIATO,
    PONTO_BEQ => W_PONTO_BEQ,
    PONTO_MUX_RT_RD => W_PONTO_MUX_RT_RD,
    PONTO_MUX_ALU_RAM => W_PONTO_MUX_ALU_RAM,
    PONTO_MUX_JMP => W_PONTO_MUX_JMP
  );

  W_CLK <= NOT W_CLK AFTER PERIODO / 2;

  main : PROCESS
  BEGIN
    W_PONTO_ESCREVE_C <= '1';
    W_PONTO_HAB_RAM <= '1';
    W_PONTO_HAB_READ <= '1';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '1';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO / 2;

    W_PONTO_ESCREVE_C <= '0';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '1';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '0';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO * 2;

    W_PONTO_ESCREVE_C <= '0';
    W_PONTO_HAB_RAM <= '1';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '1';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '1';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO;

    W_PONTO_ESCREVE_C <= '1';
    W_PONTO_HAB_RAM <= '1';
    W_PONTO_HAB_READ <= '1';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '1';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO;

    W_PONTO_ESCREVE_C <= '0';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '1';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '0';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO;

    W_PONTO_ESCREVE_C <= '1';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '1';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '0';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO * 2;

    W_PONTO_ESCREVE_C <= '0';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '0';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '1';
    WAIT FOR PERIODO;

    W_PONTO_ESCREVE_C <= '1';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '1';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '0';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO * 2;

    W_PONTO_ESCREVE_C <= '0';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '0';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '1';
    W_PONTO_OPERACAO <= '0';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '1';
    WAIT FOR PERIODO;

    W_PONTO_ESCREVE_C <= '1';
    W_PONTO_HAB_RAM <= '0';
    W_PONTO_HAB_READ <= '0';
    W_PONTO_MUX_RT_RD <= '1';
    W_PONTO_BEQ <= '0';
    W_PONTO_MUX_RT_IMEDIATO <= '0';
    W_PONTO_MUX_ALU_RAM <= '0';
    W_PONTO_OPERACAO <= '1';
    W_PONTO_HAB_WRITE <= '0';
    W_PONTO_MUX_JMP <= '0';
    WAIT FOR PERIODO;

    WAIT;
  END PROCESS main;
END test;