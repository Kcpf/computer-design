LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY RegisterFile_tb IS
END RegisterFile_tb;

ARCHITECTURE test OF RegisterFile_tb IS
  COMPONENT RegisterFile
    PORT (
      CLK : IN STD_LOGIC;
      REG_A_SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
      REG_B_SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
      REG_WRITE_SEL : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
      INPUT_DATA : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
      WRITE_ENABLE : IN STD_LOGIC := '0';
      OUT_A : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
      OUT_B : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0')
    );
  END COMPONENT;

  SIGNAL W_CLK : STD_LOGIC := '0';
  SIGNAL W_REG_A_SEL : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
  SIGNAL W_REG_B_SEL : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
  SIGNAL W_REG_WRITE_SEL : STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
  SIGNAL W_INPUT_DATA : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
  SIGNAL W_WRITE_ENABLE : STD_LOGIC := '0';
  SIGNAL W_OUT_A : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
  SIGNAL W_OUT_B : STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');

  CONSTANT PERIOD : TIME := 10 ps;

BEGIN

  RF : RegisterFile
  PORT MAP(
    CLK => W_CLK,
    REG_A_SEL => W_REG_A_SEL,
    REG_B_SEL => W_REG_B_SEL,
    REG_WRITE_SEL => W_REG_WRITE_SEL,
    INPUT_DATA => W_INPUT_DATA,
    WRITE_ENABLE => W_WRITE_ENABLE,
    OUT_A => W_OUT_A,
    OUT_B => W_OUT_B
  );

  W_CLK <= NOT W_CLK AFTER PERIOD / 2;

  main : PROCESS
  BEGIN
    W_REG_A_SEL <= "00001";
    W_REG_B_SEL <= "00010";
    W_REG_WRITE_SEL <= "00011";
    W_INPUT_DATA <= "00000000000000000000000000000001";
    W_WRITE_ENABLE <= '1';
    WAIT FOR PERIOD;
    ASSERT (W_OUT_A = "00000000000000000000000000000000") REPORT "Failure A" SEVERITY FAILURE;
    ASSERT (W_OUT_B = "00000000000000000000000000000000") REPORT "Failure B" SEVERITY FAILURE;

    W_REG_A_SEL <= "00011";
    W_REG_B_SEL <= "00011";
    W_REG_WRITE_SEL <= "00011";
    W_INPUT_DATA <= "00000000000000000000000000000001";
    W_WRITE_ENABLE <= '0';
    WAIT FOR PERIOD;
    ASSERT (W_OUT_A = "00000000000000000000000000000001") REPORT "Failure C" SEVERITY FAILURE;

    W_REG_A_SEL <= "00001";
    W_REG_B_SEL <= "00011";
    W_REG_WRITE_SEL <= "00000";
    W_INPUT_DATA <= "00000000000000000000000000000001";
    W_WRITE_ENABLE <= '1';
    WAIT FOR PERIOD;

    W_REG_A_SEL <= "00000";
    W_REG_B_SEL <= "00011";
    W_REG_WRITE_SEL <= "00001";
    W_INPUT_DATA <= "00000000000000000000000000000001";
    W_WRITE_ENABLE <= '0';
    WAIT FOR PERIOD;
    ASSERT (W_OUT_A = "00000000000000000000000000000000") REPORT "Failure D " & to_string(W_OUT_A) SEVERITY FAILURE;
  END PROCESS;
END test;