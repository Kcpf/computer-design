LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY CPU_tb IS
END CPU_tb;

ARCHITECTURE test OF CPU_tb IS
  COMPONENT CPU
    PORT (
      CLOCK_50 : IN STD_LOGIC := '0'
    );
  END COMPONENT;

  SIGNAL W_CLK : STD_LOGIC := '0';

  CONSTANT PERIODO : TIME := 10 ps;

BEGIN

  TL : CPU
  PORT MAP(
    CLOCK_50 => W_CLK
  );

  W_CLK <= NOT W_CLK AFTER PERIODO / 2;

END test;