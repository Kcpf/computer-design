LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY decoderGeneric IS
  PORT (
    entrada : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    saida : OUT STD_LOGIC_VECTOR(5 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE comportamento OF decoderGeneric IS

  CONSTANT NOP : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0000";
  CONSTANT LDA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0001";
  CONSTANT SOMA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0010";
  CONSTANT SUB : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0011";
  CONSTANT LDI : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0100";
  CONSTANT STA : STD_LOGIC_VECTOR(3 DOWNTO 0) := "0101";

BEGIN
  saida <=
    "000000" WHEN entrada = NOP ELSE
    "011010" WHEN entrada = LDA ELSE
    "010010" WHEN entrada = SOMA ELSE
    "010110" WHEN entrada = SUB ELSE
    "111000" WHEN entrada = LDI ELSE
    "001001" WHEN entrada = STA ELSE
    "000000";
END ARCHITECTURE;