LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY InstructionDecoder IS
  PORT (
    entrada : IN STD_LOGIC_VECTOR(4 DOWNTO 0) := (OTHERS => '0');
    entrada_flag_zero : IN STD_LOGIC := '0';
    entrada_flag_greater : IN STD_LOGIC := '0';
    entrada_flag_lesser : IN STD_LOGIC := '0';
    saida : OUT STD_LOGIC_VECTOR(14 DOWNTO 0) := (OTHERS => '0')
  );
END ENTITY;

ARCHITECTURE comportamento OF InstructionDecoder IS

  CONSTANT NOP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00000";
  CONSTANT LDA : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00001";
  CONSTANT SOMA : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00010";
  CONSTANT SUB : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00011";
  CONSTANT LDI : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00100";
  CONSTANT STA : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00101";
  CONSTANT JMP : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00110";
  CONSTANT JEQ : STD_LOGIC_VECTOR(4 DOWNTO 0) := "00111";
  CONSTANT CEQ : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01000";
  CONSTANT JSR : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01001";
  CONSTANT RET : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01010";
  CONSTANT CLT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01011";
  CONSTANT CGT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01100";
  CONSTANT JLT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01101";
  CONSTANT JGT : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01110";
  CONSTANT MODL : STD_LOGIC_VECTOR(4 DOWNTO 0) := "01111";
  CONSTANT DIV : STD_LOGIC_VECTOR(4 DOWNTO 0) := "10000";

  -- 14 Hab Flag Less Than
  -- 13 Hab Flag Greater Than
  -- 12 Hab escrita retorno
  -- 11 JMP
  -- 10 RET
  -- 9 JSR
  -- 8 JEQ
  -- 7 Sel MUX
  -- 6 Hab A
  -- 5, 4 e 3 Operancao
  -- 2 Hab Flag Zero
  -- 1 RD
  -- 0 WR

BEGIN
  saida <=
    "000000000000000" WHEN entrada = NOP ELSE
    "000000001010010" WHEN entrada = LDA ELSE
    "000000001000010" WHEN entrada = SOMA ELSE
    "000000001001010" WHEN entrada = SUB ELSE
    "000000011010000" WHEN entrada = LDI ELSE
    "000000000010001" WHEN entrada = STA ELSE
    "000100000000000" WHEN entrada = JMP ELSE
    "000000100000000" WHEN (entrada = JEQ AND entrada_flag_zero = '1') ELSE
    "000000000001110" WHEN entrada = CEQ ELSE
    "001001000000000" WHEN entrada = JSR ELSE
    "000010000000000" WHEN entrada = RET ELSE
    "100000000001010" WHEN entrada = CLT ELSE
    "010000000001010" WHEN entrada = CGT ELSE
    "000000100000000" WHEN (entrada = JLT AND entrada_flag_lesser = '1') ELSE
    "000000001100010" WHEN entrada = MODL ELSE
    "000000001101010" WHEN entrada = DIV ELSE
    "000000000000000"; -- NOP para os entradas Indefinidas

END ARCHITECTURE;