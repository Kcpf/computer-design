LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

ENTITY IOAddressDecoder IS
  PORT (
    ENTRADA : IN STD_LOGIC_VECTOR(8 DOWNTO 0) := (OTHERS => '0');
    RD : IN STD_LOGIC := '0';
    WR : IN STD_LOGIC := '0';
    SAIDA_RAM : OUT STD_LOGIC := '0';
    SAIDA_LED_1 : OUT STD_LOGIC := '0';
    SAIDA_LED_2 : OUT STD_LOGIC := '0';
    SAIDA_LED_FITA : OUT STD_LOGIC := '0';
    SAIDA_HEX : OUT STD_LOGIC_VECTOR(5 DOWNTO 0) := (OTHERS => '0');
    SAIDA_SW_9 : OUT STD_LOGIC := '0';
    SAIDA_SW_8 : OUT STD_LOGIC := '0';
    SAIDA_SW_7_0 : OUT STD_LOGIC := '0';
    SAIDA_KEY_3_0 : OUT STD_LOGIC_VECTOR(3 DOWNTO 0) := (OTHERS => '0');
    SAIDA_KEY_RESET : OUT STD_LOGIC := '0';
    SAIDA_CLOCK : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_0 : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_1 : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_2 : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_3 : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_RESET : OUT STD_LOGIC := '0';
    SAIDA_LIMPA_CLOCK : OUT STD_LOGIC := '0'
  );
END ENTITY;

ARCHITECTURE arch OF IOAddressDecoder IS

  COMPONENT Decoder3x8
    PORT (
      entrada : IN STD_LOGIC_VECTOR(2 DOWNTO 0);
      saida : OUT STD_LOGIC_VECTOR(7 DOWNTO 0)
    );
  END COMPONENT;

  -- DECODER BLOCO (COMPONENTE)
  SIGNAL DECODER_BLOCO_IN : STD_LOGIC_VECTOR(2 DOWNTO 0);
  SIGNAL DECODER_BLOCO_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);

  -- DECODER ENDERECO
  SIGNAL DECODER_ENDERECO_IN : STD_LOGIC_VECTOR(2 DOWNTO 0);
  SIGNAL DECODER_ENDERECO_OUT : STD_LOGIC_VECTOR(7 DOWNTO 0);

BEGIN
  DECODER_BLOCO : Decoder3x8
  PORT MAP(
    entrada => DECODER_BLOCO_IN,
    saida => DECODER_BLOCO_OUT
  );

  DECODER_ENDERECO : Decoder3x8
  PORT MAP(
    entrada => DECODER_ENDERECO_IN,
    saida => DECODER_ENDERECO_OUT
  );

  DECODER_BLOCO_IN <= ENTRADA(8 DOWNTO 6);
  DECODER_ENDERECO_IN <= ENTRADA(2 DOWNTO 0);

  SAIDA_RAM <= DECODER_BLOCO_OUT(0);

  SAIDA_LED_1 <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(4) AND
    DECODER_ENDERECO_OUT(2) AND
    WR;

  SAIDA_LED_2 <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(4) AND
    DECODER_ENDERECO_OUT(1) AND
    WR;

  SAIDA_LED_FITA <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(4) AND
    DECODER_ENDERECO_OUT(0) AND
    WR;

  SAIDA_HEX(0) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(0) AND
  WR;

  SAIDA_HEX(1) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(1) AND
  WR;

  SAIDA_HEX(2) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(2) AND
  WR;

  SAIDA_HEX(3) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(3) AND
  WR;

  SAIDA_HEX(4) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(4) AND
  WR;

  SAIDA_HEX(5) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(4) AND
  DECODER_ENDERECO_OUT(5) AND
  WR;

  SAIDA_SW_9 <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(5) AND
    DECODER_ENDERECO_OUT(2) AND
    RD;

  SAIDA_SW_8 <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(5) AND
    DECODER_ENDERECO_OUT(1) AND
    RD;

  SAIDA_SW_7_0 <= NOT(ENTRADA(5)) AND
    DECODER_BLOCO_OUT(5) AND
    DECODER_ENDERECO_OUT(0) AND
    RD;

  SAIDA_KEY_3_0(0) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(5) AND
  DECODER_ENDERECO_OUT(0) AND
  RD;

  SAIDA_KEY_3_0(1) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(5) AND
  DECODER_ENDERECO_OUT(1) AND
  RD;

  SAIDA_KEY_3_0(2) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(5) AND
  DECODER_ENDERECO_OUT(2) AND
  RD;

  SAIDA_KEY_3_0(3) <= ENTRADA(5) AND
  DECODER_BLOCO_OUT(5) AND
  DECODER_ENDERECO_OUT(3) AND
  RD;

  SAIDA_KEY_RESET <= ENTRADA(5) AND
    DECODER_BLOCO_OUT(5) AND
    DECODER_ENDERECO_OUT(4) AND
    RD;

  SAIDA_CLOCK <= ENTRADA(5) AND
    DECODER_BLOCO_OUT(5) AND
    DECODER_ENDERECO_OUT(5) AND
    RD;

  -- 511
  SAIDA_LIMPA_0 <= ENTRADA(0) AND
    ENTRADA(1) AND
    ENTRADA(2) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    ENTRADA(6) AND
    ENTRADA(7) AND
    ENTRADA(8) AND
    WR;

  -- 510
  SAIDA_LIMPA_1 <= ENTRADA(0) AND
    ENTRADA(1) AND
    ENTRADA(2) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    ENTRADA(6) AND
    ENTRADA(7) AND
    NOT(ENTRADA(8)) AND
    WR;

  -- 509
  SAIDA_LIMPA_2 <= ENTRADA(0) AND
    ENTRADA(1) AND
    ENTRADA(2) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    ENTRADA(6) AND
    NOT(ENTRADA(7)) AND
    ENTRADA(8) AND
    WR;

  -- 508
  SAIDA_LIMPA_3 <= ENTRADA(0) AND
    ENTRADA(1) AND
    ENTRADA(2) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    ENTRADA(6) AND
    NOT(ENTRADA(7)) AND
    NOT(ENTRADA(8)) AND
    WR;

  --507
  SAIDA_LIMPA_RESET <= ENTRADA(0) AND
    ENTRADA(1) AND
    ENTRADA(2) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    NOT(ENTRADA(6)) AND
    ENTRADA(7) AND
    ENTRADA(8) AND
    WR;

  -- 506
  SAIDA_LIMPA_CLOCK <= NOT(ENTRADA(0)) AND
    ENTRADA(1) AND
    NOT(ENTRADA(2)) AND
    ENTRADA(3) AND
    ENTRADA(4) AND
    ENTRADA(5) AND
    ENTRADA(6) AND
    ENTRADA(7) AND
    ENTRADA(8) AND
    WR;

END ARCHITECTURE;