LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL; --Soma (esta biblioteca =ieee)

ENTITY MainDecoder IS
  PORT (
    INSTRUCTION : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    CONTROL_WORD : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
    CONTROL_ULA : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE arch OF MainDecoder IS
  COMPONENT ControlUnit
    PORT (
      OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      CONTROL_WORD : OUT STD_LOGIC_VECTOR(8 DOWNTO 0);
      TYPE_R : OUT STD_LOGIC
    );
  END COMPONENT;

  COMPONENT DecoderFunctALU
    PORT (
      FUNCT : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      ULA_CTRL : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
  END COMPONENT;

  COMPONENT DecoderOpcodeALU
    PORT (
      OPCODE : IN STD_LOGIC_VECTOR(5 DOWNTO 0);
      ULA_CTRL : OUT STD_LOGIC_VECTOR(3 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL TYPE_R : STD_LOGIC;
  SIGNAL ULA_CTRL_FUNCT : STD_LOGIC_VECTOR(3 DOWNTO 0);
  SIGNAL ULA_CTRL_OPCODE : STD_LOGIC_VECTOR(3 DOWNTO 0);

BEGIN
  ControlUnit_PORT_MAP : ControlUnit
  PORT MAP(
    OPCODE => INSTRUCTION(31 DOWNTO 26),
    CONTROL_WORD => CONTROL_WORD,
    TYPE_R => TYPE_R
  );

  DecoderFunctALU_PORT_MAP : DecoderFunctALU
  PORT MAP(
    FUNCT => INSTRUCTION(5 DOWNTO 0),
    ULA_CTRL => ULA_CTRL_FUNCT
  );

  DecoderOpcodeALU_PORT_MAP : DecoderOpcodeALU
  PORT MAP(
    OPCODE => INSTRUCTION(31 DOWNTO 26),
    ULA_CTRL => ULA_CTRL_OPCODE
  );

  CONTROL_ULA <= ULA_CTRL_OPCODE WHEN TYPE_R = '0' ELSE
    ULA_CTRL_FUNCT;

END ARCHITECTURE;