LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL; -- Biblioteca IEEE para funções aritméticas

ENTITY ALU IS
  PORT (
    INPUT_A : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
    INPUT_B : IN STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
    SEL : IN STD_LOGIC := '0';
    OUTPUT : OUT STD_LOGIC_VECTOR(31 DOWNTO 0) := (OTHERS => '0');
    FLAG_EQUAL : OUT STD_LOGIC := '0'
  );
END ENTITY;

ARCHITECTURE arch OF ALU IS
  SIGNAL SUM : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL SUB : STD_LOGIC_VECTOR(31 DOWNTO 0);

BEGIN
  SUM <= STD_LOGIC_VECTOR(unsigned(INPUT_A) + unsigned(INPUT_B));
  SUB <= STD_LOGIC_VECTOR(unsigned(INPUT_A) - unsigned(INPUT_B));

  OUTPUT <= SUM WHEN (SEL = '1') ELSE
    SUB;
  FLAG_EQUAL <= '1' WHEN (INPUT_A = INPUT_B) ELSE
    '0';
END ARCHITECTURE;