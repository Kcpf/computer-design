LIBRARY IEEE;
USE IEEE.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

ENTITY ROM IS
  GENERIC (
    dataWidth : NATURAL := 4;
    addrWidth : NATURAL := 3
  );
  PORT (
    Endereco : IN STD_LOGIC_VECTOR (addrWidth - 1 DOWNTO 0) := (OTHERS => '0');
    Dado : OUT STD_LOGIC_VECTOR (dataWidth - 1 DOWNTO 0) := (OTHERS => '0')
  );
END ENTITY;

ARCHITECTURE assincrona OF ROM IS

  TYPE blocoMemoria IS ARRAY(0 TO 2 ** addrWidth - 1) OF STD_LOGIC_VECTOR(dataWidth - 1 DOWNTO 0);

  FUNCTION initMemory
    RETURN blocoMemoria IS VARIABLE tmp : blocoMemoria := (OTHERS => (OTHERS => '0'));
  BEGIN

    -- SETUP:
    tmp(0) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(1) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(2) := "00101" & "00" & "100000001"; -- STA %R0, @257
    tmp(3) := "00101" & "00" & "100000010"; -- STA %R0, @258
    tmp(4) := "00101" & "00" & "100100000"; -- STA %R0, @288
    tmp(5) := "00101" & "00" & "100100001"; -- STA %R0, @289
    tmp(6) := "00101" & "00" & "100100010"; -- STA %R0, @290
    tmp(7) := "00101" & "00" & "100100011"; -- STA %R0, @291
    tmp(8) := "00101" & "00" & "100100100"; -- STA %R0, @292
    tmp(9) := "00101" & "00" & "100100101"; -- STA %R0, @293
    tmp(10) := "00101" & "00" & "000000000"; -- STA %R0, @0
    tmp(11) := "00101" & "00" & "000000110"; -- STA %R0, @6
    tmp(12) := "00101" & "00" & "000000111"; -- STA %R0, @7
    tmp(13) := "00101" & "00" & "000001000"; -- STA %R0, @8
    tmp(14) := "00101" & "00" & "000001001"; -- STA %R0, @9
    tmp(15) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(16) := "00101" & "00" & "000001011"; -- STA %R0, @11
    tmp(17) := "00101" & "00" & "000001100"; -- STA %R0, @12
    tmp(18) := "00100" & "00" & "000000001"; -- LDI %R0, $1
    tmp(19) := "00101" & "00" & "000000001"; -- STA %R0, @1
    tmp(20) := "00100" & "00" & "000000010"; -- LDI %R0, $2
    tmp(21) := "00101" & "00" & "000000010"; -- STA %R0, @2
    tmp(22) := "00100" & "00" & "000000100"; -- LDI %R0, $4
    tmp(23) := "00101" & "00" & "000000011"; -- STA %R0, $3
    tmp(24) := "00100" & "00" & "000000110"; -- LDI %R0, $6
    tmp(25) := "00101" & "00" & "000000100"; -- STA %R0, $4
    tmp(26) := "00100" & "00" & "000001010"; -- LDI %R0, $10
    tmp(27) := "00101" & "00" & "000000101"; -- STA %R0, $5
    tmp(28) := "01001" & "00" & "010001110"; -- JSR @CONFIGURA_RELOGIO

    -- LOOP:
    tmp(29) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(30) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(31) := "00111" & "00" & "000100001"; -- JEQ @VERIFICA_FLAG_RAPIDO
    tmp(32) := "01001" & "00" & "010001110"; -- JSR @CONFIGURA_RELOGIO

    -- VERIFICA_FLAG_RAPIDO:
    tmp(33) := "00001" & "00" & "101100000"; -- LDA %R0, @352
    tmp(34) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(35) := "00111" & "00" & "000100101"; -- JEQ @INICIO_LOOP
    tmp(36) := "01001" & "00" & "010000011"; -- JSR @TROCA_BASE

    -- INICIO_LOOP:
    tmp(37) := "00001" & "00" & "000001100"; -- LDA %R0, @12
    tmp(38) := "01000" & "00" & "000000001"; -- CEQ %R0, @1
    tmp(39) := "00111" & "00" & "000101101"; -- JEQ @SAMPA
    tmp(40) := "00001" & "00" & "101100101"; -- LDA %R0, @357
    tmp(41) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(42) := "00111" & "00" & "000110001"; -- JEQ @DISPLAY
    tmp(43) := "01001" & "00" & "000111110"; -- JSR @INCREMENTO
    tmp(44) := "00110" & "00" & "000110001"; -- JMP @DISPLAY

    -- SAMPA:
    tmp(45) := "00001" & "00" & "101100110"; -- LDA %R0, @358
    tmp(46) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(47) := "00111" & "00" & "000110001"; -- JEQ @DISPLAY
    tmp(48) := "01001" & "00" & "000111110"; -- JSR @INCREMENTO

    -- DISPLAY:
    tmp(49) := "00001" & "00" & "000000110"; -- LDA %R0, @6
    tmp(50) := "00101" & "00" & "100100000"; -- STA %R0, @288
    tmp(51) := "00001" & "01" & "000000111"; -- LDA %R1, @7
    tmp(52) := "00101" & "01" & "100100001"; -- STA %R1, @289
    tmp(53) := "00001" & "00" & "000001000"; -- LDA %R0, @8
    tmp(54) := "00101" & "00" & "100100010"; -- STA %R0, @290
    tmp(55) := "00001" & "01" & "000001001"; -- LDA %R1, @9
    tmp(56) := "00101" & "01" & "100100011"; -- STA %R1, @291
    tmp(57) := "00001" & "00" & "000001010"; -- LDA %R0, @10
    tmp(58) := "00101" & "00" & "100100100"; -- STA %R0, @292
    tmp(59) := "00001" & "01" & "000001011"; -- LDA %R1, @11
    tmp(60) := "00101" & "01" & "100100101"; -- STA %R1, @293
    tmp(61) := "00110" & "00" & "000011101"; -- JMP @LOOP

    -- INCREMENTO:
    tmp(62) := "00001" & "00" & "000001100"; -- LDA %R0, @12
    tmp(63) := "01000" & "00" & "000000001"; -- CEQ %R0, @1
    tmp(64) := "00111" & "00" & "001000100"; -- JEQ @SAMPA2
    tmp(65) := "00100" & "00" & "000000001"; -- LDI %R0, $1
    tmp(66) := "00101" & "00" & "111111010"; -- STA %R0, @506
    tmp(67) := "00110" & "00" & "001000110"; -- JMP @INCREMENTO_INICIO

    -- SAMPA2:
    tmp(68) := "00100" & "00" & "000000001"; -- LDI %R0, $1
    tmp(69) := "00101" & "00" & "111111001"; -- STA %R0, @505

    -- INCREMENTO_INICIO:
    tmp(70) := "00001" & "00" & "000000110"; -- LDA %R0, @6
    tmp(71) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(72) := "01000" & "00" & "000000101"; -- CEQ %R0, @5
    tmp(73) := "00111" & "00" & "001001100"; -- JEQ @INCREMENTA_SEGUNDO_DEC
    tmp(74) := "00101" & "00" & "000000110"; -- STA %R0, @6
    tmp(75) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTA_SEGUNDO_DEC:
    tmp(76) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(77) := "00101" & "00" & "000000110"; -- STA %R0, @6
    tmp(78) := "00001" & "00" & "000000111"; -- LDA %R0, @7
    tmp(79) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(80) := "01000" & "00" & "000000100"; -- CEQ %R0, @4
    tmp(81) := "00111" & "00" & "001010100"; -- JEQ @INCREMENTA_MINUTO
    tmp(82) := "00101" & "00" & "000000111"; -- STA %R0, @7
    tmp(83) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTA_MINUTO:
    tmp(84) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(85) := "00101" & "00" & "000000111"; -- STA %R0, @7
    tmp(86) := "00001" & "00" & "000001000"; -- LDA %R0, @8
    tmp(87) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(88) := "01000" & "00" & "000000101"; -- CEQ %R0, @5
    tmp(89) := "00111" & "00" & "001011100"; -- JEQ @INCREMENTA_MINUTO_DEC
    tmp(90) := "00101" & "00" & "000001000"; -- STA %R0, @8
    tmp(91) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTA_MINUTO_DEC:
    tmp(92) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(93) := "00101" & "00" & "000001000"; -- STA %R0, @8
    tmp(94) := "00001" & "00" & "000001001"; -- LDA %R0, @9
    tmp(95) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(96) := "01000" & "00" & "000000100"; -- CEQ %R0, @4
    tmp(97) := "00111" & "00" & "001100100"; -- JEQ @INCREMENTA_HORA
    tmp(98) := "00101" & "00" & "000001001"; -- STA %R0, @9
    tmp(99) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTA_HORA:
    tmp(100) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(101) := "00101" & "00" & "000001001"; -- STA %R0, @9
    tmp(102) := "00001" & "00" & "000001011"; -- LDA %R0, @11
    tmp(103) := "01000" & "00" & "000000010"; -- CEQ %R0, @2
    tmp(104) := "00111" & "00" & "001110101"; -- JEQ @INCREMENTO_OVERFLOW
    tmp(105) := "00001" & "00" & "000001010"; -- LDA %R0, @10
    tmp(106) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(107) := "01000" & "00" & "000000101"; -- CEQ %R0, @5
    tmp(108) := "00111" & "00" & "001101111"; -- JEQ @INCREMENTO_HORA_DEC
    tmp(109) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(110) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTO_HORA_DEC:
    tmp(111) := "00100" & "00" & "000000000"; -- LDI %R0, $0
    tmp(112) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(113) := "00001" & "00" & "000001011"; -- LDA %R0, @11
    tmp(114) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(115) := "00101" & "00" & "000001011"; -- STA %R0, @11
    tmp(116) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTO_OVERFLOW:
    tmp(117) := "00001" & "00" & "000001010"; -- LDA %R0, $10
    tmp(118) := "00010" & "00" & "000000001"; -- SOMA %R0, @1
    tmp(119) := "01000" & "00" & "000000011"; -- CEQ %R0, @3
    tmp(120) := "00111" & "00" & "001111011"; -- JEQ @INCREMENTO_RESET
    tmp(121) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(122) := "01010" & "00" & "000000000"; -- RET

    -- INCREMENTO_RESET:
    tmp(123) := "00001" & "00" & "000000000"; -- LDA %R0, @0
    tmp(124) := "00101" & "00" & "000000110"; -- STA %R0, @6
    tmp(125) := "00101" & "00" & "000000111"; -- STA %R0, @7
    tmp(126) := "00101" & "00" & "000001000"; -- STA %R0, @8
    tmp(127) := "00101" & "00" & "000001001"; -- STA %R0, @9
    tmp(128) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(129) := "00101" & "00" & "000001011"; -- STA %R0, @11
    tmp(130) := "01010" & "00" & "000000000"; -- RET

    -- TROCA_BASE:
    tmp(131) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(132) := "00101" & "00" & "111111111"; -- STA %R0, @511
    tmp(133) := "00001" & "00" & "000001100"; -- LDA %R0, @12
    tmp(134) := "01000" & "00" & "000000001"; -- CEQ %R0, @1
    tmp(135) := "00111" & "00" & "010001011"; -- JEQ @VIRA_0
    tmp(136) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(137) := "00101" & "00" & "000001100"; -- STA %R0, @12
    tmp(138) := "01010" & "00" & "000000000"; -- RET

    -- VIRA_0:
    tmp(139) := "00001" & "00" & "000000000"; -- LDA %R0, @0
    tmp(140) := "00101" & "00" & "000001100"; -- STA %R0, @12
    tmp(141) := "01010" & "00" & "000000000"; -- RET

    -- CONFIGURA_RELOGIO:
    tmp(142) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(143) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_SEG_UNI:
    tmp(144) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(145) := "00101" & "00" & "000000110"; -- STA %R0, @6
    tmp(146) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(147) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(148) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(149) := "00111" & "00" & "010010000"; -- JEQ @CONFIGURA_SEG_UNI
    tmp(150) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(151) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_RELOGIO_SEG_DEC:
    tmp(152) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(153) := "00101" & "00" & "000000111"; -- STA %R0, @7
    tmp(154) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(155) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(156) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(157) := "00111" & "00" & "010011000"; -- JEQ @CONFIGURA_RELOGIO_SEG_DEC
    tmp(158) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(159) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_RELOGIO_MIN_UNI:
    tmp(160) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(161) := "00101" & "00" & "000001000"; -- STA %R0, @8
    tmp(162) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(163) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(164) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(165) := "00111" & "00" & "010100000"; -- JEQ @CONFIGURA_RELOGIO_MIN_UNI
    tmp(166) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(167) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_RELOGIO_MIN_DEC:
    tmp(168) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(169) := "00101" & "00" & "000001001"; -- STA %R0, @9
    tmp(170) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(171) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(172) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(173) := "00111" & "00" & "010101000"; -- JEQ @CONFIGURA_RELOGIO_MIN_DEC
    tmp(174) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(175) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_RELOGIO_HORA_UNI:
    tmp(176) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(177) := "00101" & "00" & "000001010"; -- STA %R0, @10
    tmp(178) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(179) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(180) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(181) := "00111" & "00" & "010110000"; -- JEQ @CONFIGURA_RELOGIO_HORA_UNI
    tmp(182) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(183) := "00101" & "00" & "111111110"; -- STA %R0, @510

    -- CONFIGURA_RELOGIO_HORA_DEC:
    tmp(184) := "00001" & "00" & "101000000"; -- LDA %R0, @320
    tmp(185) := "00101" & "00" & "000001011"; -- STA %R0, @11
    tmp(186) := "00101" & "00" & "100000000"; -- STA %R0, @256
    tmp(187) := "00001" & "00" & "101100001"; -- LDA %R0, @353
    tmp(188) := "01000" & "00" & "000000000"; -- CEQ %R0, @0
    tmp(189) := "00111" & "00" & "010111000"; -- JEQ @CONFIGURA_RELOGIO_HORA_DEC
    tmp(190) := "00001" & "00" & "000000001"; -- LDA %R0, @1
    tmp(191) := "00101" & "00" & "111111110"; -- STA %R0, @510
    tmp(192) := "01010" & "00" & "000000000"; -- RET

    RETURN tmp;
  END initMemory;

  SIGNAL memROM : blocoMemoria := initMemory;

BEGIN
  Dado <= memROM (to_integer(unsigned(Endereco)));
END ARCHITECTURE;